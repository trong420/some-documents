module top1;
  logic clk, enb, reset_n;
  logic [2:0] req, ack, done, intrpt;
    
 m_equivalent dut(.*);
 
       default clocking @(posedge clk); endclocking
    
    
endmodule : top1
//
