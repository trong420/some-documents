module top1;
logic clk, a, b;
     
 x dut(.*);
 
       default clocking @(posedge clk); endclocking
      
endmodule : top1
//
