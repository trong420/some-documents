module top1;
    logic clk, bus_select, bus1, req1, ack1, req2, ack2;
  if_else_prop dut (.*);
     
    default clocking cb_clk @ (clk);
    endclocking 
  endmodule : top1
